module main

import io

fn main() {
}