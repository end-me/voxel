module main

import server

fn main() {
	server.new(4089)
}