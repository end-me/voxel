module packets

enum State {
	Handshake
	Status
	Login
	Play
}